library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity rq_ctrl is
    Port (
    );
end rq_ctrl;

architecture Behavioral of rq_ctrl is

end Behavioral;