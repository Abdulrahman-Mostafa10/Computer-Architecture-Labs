LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY mv_ctrl IS
    PORT (
    );
END mv_ctrl;

ARCHITECTURE Behavioral OF mv_ctrl IS

END Behavioral;