LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY rq_ctrl IS
    PORT (
    );
END rq_ctrl;

ARCHITECTURE Behavioral OF rq_ctrl IS

END Behavioral;