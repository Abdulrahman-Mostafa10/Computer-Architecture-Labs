library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity elevator_tb is
end elevator_tb;

architecture Behavioral of elevator_tb is

end Behavioral;