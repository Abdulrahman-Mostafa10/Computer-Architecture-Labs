LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY elevator IS
    PORT (
    );
END elevator;

ARCHITECTURE Behavioral OF elevator IS

END Behavioral;