library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity mv_ctrl is
    Port (
    );
end mv_ctrl;

architecture Behavioral of mv_ctrl is

end Behavioral;