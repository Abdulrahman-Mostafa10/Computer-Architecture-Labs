library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity elevator is
    Port (
    );
end elevator;

architecture Behavioral of elevator is

end Behavioral;